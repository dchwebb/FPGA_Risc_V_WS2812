.SysClk_Rst_GenMon_inst.set_clk_freq_mhz(50);
.SysClk_Rst_GenMon_inst.start_clk();
